`timescale 1ns / 1ps
module _tb;
    parameter real FREQ  = 300.0            ; // MHZ
    parameter real CYCLE = 1.0 * 1000.0/FREQ;

    /*------------------------------------------------------------------------------
    --   Signals declaration
    ------------------------------------------------------------------------------*/



    /*------------------------------------------------------------------------------
    --  DUT
    ------------------------------------------------------------------------------*/



    /*------------------------------------------------------------------------------
    --  TASKS
    ------------------------------------------------------------------------------*/
    task automatic cycles(input int number, ref bit clk,input real time_cycle);
        repeat (number) @(posedge clk) #(time_cycle/10.0);
    endtask : cycles


    /*------------------------------------------------------------------------------
    --   Behavior
    ------------------------------------------------------------------------------*/
    always #(CYCLE/2.0) clk_ = !clk_  ;

    initial begin
        rst = 1;
        cycles(5,clk_,CYCLE);
        rst = 0;
        cycles(5,clk_,CYCLE);

    end
endmodule
